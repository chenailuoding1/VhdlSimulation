library IEEE;

use IEEE.STD_LOGIC_1164.ALL;

use IEEE.std_logic_unsigned.All;

USE ieee.numeric_std.ALL;

--指令（instruction）统一为std_logic数据类型，值（value，signal）统一为STD_LOGIC_VECTOR ( 31 downto 0 )数据类型
entity IT is
port(
	in_32IT_32IT_32ms_inte_time_star_inst:in STD_LOGIC_VECTOR ( 31 downto 0 )--in_32ITI_32IT_32ms interrupt timer start instruction
);
end IT;
architecture Behavioral of IT is
begin
--需要用户补全的信息




end Behavioral;
